//incomplete
module registerAverage(
    input i_clk,
    input i_reset,
    input i_enableWrite,
    input [15:0] i_selWrite,
    input [9:0] i_data0,
    input [9:0] i_data1,
    input [9:0] i_data2,
    output [159:0] o_ave,
);
endmodule