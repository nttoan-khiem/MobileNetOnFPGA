module ramConvWrp(
    
);

endmodule